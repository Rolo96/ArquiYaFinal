library verilog;
use verilog.vl_types.all;
entity decobench is
end decobench;
