library verilog;
use verilog.vl_types.all;
entity add is
end add;
